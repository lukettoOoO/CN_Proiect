library verilog;
use verilog.vl_types.all;
entity restoring_tb is
end restoring_tb;
