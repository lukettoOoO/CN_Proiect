module smtoc2_tb;
  reg [7:0] x, y;
  wire [7:0] x_c2, y_c2;
  
  smtoc2 inst (
    .x(x),
    .y(y),
    .x_c2(x_c2),
    .y_c2(y_c2)
  );
  
  initial begin
    x = 8'b00000101; //5
    y = 8'b10000101; //-5
    #10;

    x = 8'b00000001; //1
    y = 8'b10000001; //-1
    #10;

    x = 8'b11111111; //-127
    y = 8'b01111111; //127
    #10;

    x = 8'b00000000; // 0
    y = 8'b10000000; //-128
    #10;

    x = 8'b00000010; //2 
    y = 8'b10000010; //-2
    #10;
  end
  
endmodule