library verilog;
use verilog.vl_types.all;
entity rca8_tb is
end rca8_tb;
