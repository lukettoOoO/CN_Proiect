module c2tosm_tb; 
  reg [7:0] x;
  wire [7:0] sm;
  
  c2tosm inst (
    .x(x),
    .sm(sm)
  );
  
  initial begin
    x = 8'b00000101;  //5
    #10;
    //sm = 00000101

    x = 8'b11111011;  //-5
    #10;

    x = 8'b00000000;  //0
    #10;
    //sm = 00000000

    x = 8'b01111111;  //127
    #10;
    //sm = 01111111

    x = 8'b10000001;  //-127
    #10;
    //sm = 10000001

    x = 8'b10000000;  //-128
    #10;
    //sm = 10000000
  end
  
endmodule